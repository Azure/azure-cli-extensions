61 38 6b 92 16 4b cc ac 6f d4 02 5c 6f 62 79 b9 
8e 62 ae 07 02 1c dc 73 5b 7a 51 e7 56 4e 4a b0 
54 4a 93 2e 6b dd 3c b5 8b 60 fa 80 b1 80 1b 89 
1e 4d 7d 86 8e 25 76 58 24 8d 21 87 83 06 88 d6 
a4 fd 94 9c 66 b6 db ee 92 46 f0 25 fc 84 bb f5 
3f d9 49 28 ea 54 6a 2a 33 fa e0 47 eb 22 af 91 
d4 34 a6 d9 fe 58 cb 54 03 35 d6 45 40 96 4e f3 
31 ea 78 20 45 e9 f2 3a de cb 38 53 c0 9c b2 b7 
12 9e 57 d9 f6 1b cb 20 23 8c 86 d3 40 da 84 c3 
22 5b 48 61 63 e2 5f 5f 43 6d 8f 41 fc ce c1 87 
33 e1 e2 61 63 e2 5f 5